package my_pkg;
  `include "apb_master_transaction.sv"
  `include "apb_master_generator.sv"
  `include "apb_master_driver.sv"
  `include "apb_master_monitor.sv"
  `include "apb_master_scoreboard.sv"
  `include "apb_master_environment.sv"
 // `include "apb_master_test.sv"
endpackage
